----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.12.2020 19:27:01
-- Design Name: 
-- Module Name: pwm_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.package_dsed.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pwm_tb is
end pwm_tb;

architecture Behavioral of pwm_tb is

component pwm 
    Port ( clk_12megas : in STD_LOGIC;
           reset : in STD_LOGIC;
           en_2_cycles : in STD_LOGIC;
           sample_in : in STD_LOGIC_VECTOR (sample_size-1 downto 0);
           sample_request : out STD_LOGIC;
           pwm_pulse : out STD_LOGIC);
end component;

component enables
    Port ( clk_12megas : in STD_LOGIC;
           reset : in STD_LOGIC;
           clk_3megas : out STD_LOGIC;
           en_2_cycles : out STD_LOGIC;
           en_4_cycles : out STD_LOGIC);
end component;

signal clk_12megas, reset, enable_2_cycles_aux, sample_request, pwm_pulse, clk_3megas, en_4_cycles : std_logic :='0';
signal sample_in: STD_LOGIC_VECTOR (7 downto 0):= "00000000";
constant clk_period : time := 10 ns;

begin

EN2: enables
        port map (
            clk_12megas => clk_12megas, 
            reset => reset,
            clk_3megas => clk_3megas,
            en_2_cycles => enable_2_cycles_aux, 
            en_4_cycles => en_4_cycles);

DUT: pwm 
        port map (
            clk_12megas => clk_12megas, 
            reset => reset,
            en_2_cycles => enable_2_cycles_aux,
            sample_in => sample_in,  
            sample_request => sample_request, 
            pwm_pulse => pwm_pulse);
            
clk_process :process
             begin
             clk_12megas <= '0';
             wait for clk_period/2;
                clk_12megas <= '1';
             wait for clk_period/2;
             end process;        
                 
sim_proc:   process
            begin
            reset<='1';
            wait for 100ns;
            reset<='0';
            wait for 100ns;
            sample_in<= "00000000";
            wait for 300 us;
            sample_in<= "00101001";
            wait for 300 us;
            sample_in<= "11111111";
            wait;
            end process;


end Behavioral;
