package package_dsed is
    constant sample_size: integer :=8;
end package_dsed;  